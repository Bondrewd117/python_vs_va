*================================================================
* Automated SPICE simulation for comparison
*================================================================

.control
pre_osdi /foss/designs/Capibara_tuto/MEMS/rram_v1_with_monitors.osdi
.endc

.options num_threads=8
.options method=gear
.options maxstep=2u
.options reltol=1e-4
.options abstol=1e-12

.subckt rram_v1 TE BE X_OUT G_OUT VM_OUT IS_OUT IM_OUT
N1 TE BE X_OUT G_OUT VM_OUT IS_OUT IM_OUT rram_v1_model
.ends

.model rram_v1_model rram_v1_va 
+ x0=0.0 Ron=13e3 Roff=460e3 tau=6e-5 T=108.5
+ Von_threshold=0.2 Voff=-0.1 phi=0.88
+ Af=1e-7 Ar=1e-7 Bf=8 Br=8

* Circuit
Vin V_input 0 SIN(0 0.4 10)
Rs V_input TE 10k
Xmem TE 0 X_mon G_mon Vm_mon Is_mon Im_mon rram_v1

.tran 2u 200m

.control
    save all
    run
    set wr_singlescale
    set wr_vecnames
    option numdgt=15
    wrdata /foss/designs/Capibara_tuto/MEMS/tmp/spice_results.txt time v(V_input) v(Vm_mon) v(X_mon) v(G_mon) v(Im_mon) v(Is_mon) i(Vin)
    quit
.endc

.end
